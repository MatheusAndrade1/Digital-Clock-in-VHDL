----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 23.08.2019 19:35:48
-- Design Name: 
-- Module Name: Decod - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity Decod is
  Port (e: in STD_LOGIC_VECTOR (1 downto 0);
        an: out STD_LOGIC_VECTOR (3 downto 0) );
end Decod;

architecture Behavioral of Decod is

begin

with e select
    an <= "1110" when "00",
          "1101" when "01",
          "1011" when "10",
          "0111" when "11",
          "1111" when others;

end Behavioral;
